package ahb_pkg;                       // package declaration
  
  import uvm_pkg::*; 
  `include "uvm_macros.svh"                  // import UVM package

//====================================
// Includes
//====================================
`include "interface.sv"      
`include "ahb_seq_item.sv"
`include "ahb_driver.sv"
`include "ahb_monitor.sv"
`include "ahb_agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "ahb_sequence.sv"
`include "test.sv"
  
endpackage 